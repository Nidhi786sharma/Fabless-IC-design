module parity_encoder(in,out);
output [2:0]out;
reg [2:0]out;
input [7:0]in;
wire [7:0]in;

