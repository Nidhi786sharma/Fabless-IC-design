module or_gate(out,a,b);
output out;
input a,b;
or o1(out,a,b);
endmodule
